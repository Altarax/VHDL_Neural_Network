--! Import libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package types is

    type int_array is array (natural range <>) of integer;
    
end package types;

package body types is
    
end package body types;