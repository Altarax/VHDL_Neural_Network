--! Import libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--! Import custom library
library work;
use work.types.all;

--! \brief Activation function
--! \details
entity act_funct is
    generic (

    );
    port (

    );
end entity neuron;

architecture rtl of act_func is

    
begin
    
    
end architecture rtl;