--! Import libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--! Import custom library
library work;
use work.types.all;

--! \brief Neural Network
--! \details
entity network is
    port (

    );
end entity network;

architecture rtl of network is

    
begin
    
    
end architecture rtl;