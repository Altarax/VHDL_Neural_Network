--! Import libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--! Import custom library
library work;
use work.types.all;

--! \brief Simple Neuron
--! \details
entity neuron is
	generic (
        
	);
    port (

    );
end entity neuron;

architecture rtl of neuron is

begin

    
end architecture rtl;